--main entity of the proj no. 4, DE2_mul 
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY DE2_mul IS
	PORT(SW : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		  
		  
		  HEX6: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX4: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX1: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX0: OUT STD_LOGIC_VECTOR(0 TO 6));


END DE2_mul;

ARCHITECTURE Behaviour OF DE2_mul IS
COMPONENT mul
	PORT(A,B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 P: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT hex_to_disp
    Port ( HEX_NUM : IN STD_LOGIC_VECTOR (3 downto 0);
           TO_DISP : OUT  STD_LOGIC_VECTOR (0 to 6));
END COMPONENT;

SIGNAL PRODUCT:STD_LOGIC_VECTOR(0 TO 6);
BEGIN

mul1:mul PORT MAP(SW(11 DOWNTO 8),SW(3 DOWNTO 0),PRODUCT);

disp6:hex_to_disp PORT MAP(SW(11 DOWNTO 8),HEX6);
disp4:hex_to_disp PORT MAP(SW(3 DOWNTO 0),HEX4);

disp1:hex_to_disp PORT MAP(PRODUCT(7 DOWNTO 4),HEX1);
disp0:hex_to_disp PORT MAP(PRODUCT(3 DOWNTO 0),HEX0);

END Behaviour;