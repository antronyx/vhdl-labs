LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--main code
ENTITY RCA_8bit IS
	PORT( 	 	 SW: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			KEY0,KEY1: IN STD_LOGIC; -- respectively reset and clock
			  LEDG[8]: OUT STD_LOGIC;
				  LEDR: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
				  HEX7: OUT STD_LOGIC_VECTOR(0 TO 6);
				  HEX6: OUT STD_LOGIC_VECTOR(0 TO 6);
				  HEX5: OUT STD_LOGIC_VECTOR(0 TO 6);
				  HEX4: OUT STD_LOGIC_VECTOR(0 TO 6);
				  HEX1: OUT STD_LOGIC_VECTOR(0 TO 6);
				  HEX0: OUT STD_LOGIC_VECTOR(0 TO 6)
	);

END RCA_8bit;


ARCHITECTURE Behaviour OF 8bit_RCA IS
	COMPONENT SAdd_8bit 
		PORT(A,B: IN STD_LOGIC_VECTOR(7 DOWNTO 0); 	 	 
				 S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
  C_in,CLK,RST: IN STD_LOGIC;
			C_out: OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT hex_to_disp 
	PORT (HEX_NUM: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			TO_DISP: OUT STD_LOGIC_VECTOR(0 TO 6);
			OVFL:IN STD_LOGIC);
	END COMPONENT;
	
SIGNAL RESULT : STD_LOGIC_VECTOR(7 DOWNTO 0);	
SIGNAL NUM1:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL NUM2:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL OVFL_STATUS:STD_LOGIC;
BEGIN
	
	NUM1<=SW(15 DOWNTO 8);
	NUM2<=SW(7 DOWNTO 0);
	ADD0:SAdd_8bit PORT MAP(NUM1,NUM2,RESULT,'0',KEY1,KEY0,OVFL_STATUS);
	
	--------INPUTS DISPAY-------------------------------
	hex7:hex_to_disp PORT MAP(NUM1(7 DOWNTO 4),HEX7,'0');
	hex6:hex_to_disp PORT MAP(NUM1(3 DOWNTO 0),HEX6,'0');
	
	hex5:hex_to_disp PORT MAP(NUM2(7 DOWNTO 4),HEX5,'0');
	hex4:hex_to_disp PORT MAP(NUM2(3 DOWNTO 0),HEX4,'0');
	-----------------------------------------------------
	
	-------OUTPUT DISPLAY--------------------------------
	hex1:hex_to_disp PORT MAP(RESULT(7 DOWNTO 4),HEX1,OVFL_STATUS);
	hex0:hex_to_disp PORT MAP(RESULT(3 DOWNTO 0),HEX0,OVFL_STATUS);
	LEDG[8]<=OVFL_OCCURRED;
	------------------------------------------------------
	

END Behaviour;